library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mem_fondo is
	Port(
		NIVEL : IN integer;
		FILA : IN integer;
		COLUMNA : IN integer;
		COLORES : OUT integer);	
end mem_fondo;

architecture Behavioral of mem_fondo is

type mem_matrix is array (0 to 23, 0 to 31) of integer;

constant inicio : mem_matrix := (
	(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
	(1,1,1,1,2,12,12,12,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
	(1,1,1,2,12,12,12,12,12,12,12,12,1,2,12,12,1,1,2,12,12,12,1,1,2,12,2,12,1,1,1,1),
	(1,1,1,2,12,13,15,15,15,15,15,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1),
	(1,1,1,2,12,13,15,12,12,13,15,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1),
	(1,1,1,2,12,13,15,12,12,12,12,12,12,13,15,15,12,12,13,15,15,15,12,12,13,15,13,15,12,12,12,1),
	(1,1,1,2,12,13,15,12,13,15,15,12,13,15,12,13,15,12,13,15,12,13,15,12,13,15,15,15,12,12,12,1),
	(1,1,1,2,12,13,15,12,12,13,15,12,13,15,15,15,15,12,13,15,15,15,12,12,12,13,15,12,12,12,12,1),
	(1,1,1,2,12,13,15,12,12,13,15,12,13,15,12,13,15,12,13,15,12,13,15,12,12,13,15,12,12,12,12,1),
	(1,1,1,2,12,13,15,15,15,15,15,12,13,15,12,13,15,12,13,15,12,13,15,12,12,13,15,12,12,12,1,1),
	(1,1,1,2,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1,1,1),
	(1,1,1,1,2,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1,1,1,1),
	(1,1,1,1,1,1,2,12,12,12,1,1,2,12,1,2,12,1,2,12,1,2,12,1,1,2,12,1,1,1,1,1),
	(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
	(1,1,1,1,1,2,12,12,12,12,1,2,12,12,12,1,1,2,12,1,1,2,12,12,1,1,2,12,12,12,1,1),
	(1,1,1,2,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1),
	(1,1,1,2,12,12,13,15,15,15,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1),
	(1,1,1,2,12,13,15,12,12,12,12,13,15,15,15,12,12,13,15,12,12,13,15,15,12,12,13,15,15,15,12,1),
	(1,1,1,2,12,12,13,15,15,12,12,12,13,15,12,12,13,15,12,15,12,13,15,13,15,12,12,13,15,12,12,1),
	(1,1,1,2,12,12,12,12,13,15,12,12,13,15,12,12,13,15,15,15,12,13,15,15,12,12,12,13,15,12,12,1),
	(1,1,1,2,12,13,15,15,15,12,12,12,13,15,12,12,13,15,12,15,12,13,15,13,15,12,12,13,15,12,12,1),
	(1,1,1,2,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1,1),
	(1,1,1,1,1,2,12,12,12,1,1,1,2,12,1,1,2,12,2,12,1,2,12,2,12,1,1,2,12,1,1,1),
	(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1)
	);

constant nivel_1 : mem_matrix := (
	(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
	(1,1,1,7,7,7,8,7,7,7,7,7,7,7,7,7,7,7,8,9,9,8,8,9,8,8,8,8,2,2,2,1),
	(1,1,1,7,7,7,9,7,7,8,8,9,8,8,7,7,9,8,8,9,9,8,7,7,7,7,7,8,8,2,2,1),
	(1,1,1,8,9,7,8,7,8,9,7,7,7,8,7,8,8,7,9,7,7,8,8,8,9,8,8,8,8,7,2,1),
	(1,1,1,7,7,7,7,7,8,7,7,8,7,8,7,7,7,8,8,7,7,7,7,7,7,7,7,7,7,7,7,1),
	(1,1,1,8,7,8,8,7,8,7,7,8,9,14,2,2,7,8,7,9,8,8,8,7,8,8,8,14,14,8,7,1),
	(1,1,1,7,7,7,8,7,7,7,7,7,8,14,14,8,7,7,7,7,8,8,8,7,8,2,2,14,8,14,8,1),
	(1,1,1,7,7,7,9,7,7,14,8,7,8,7,7,8,8,9,7,7,7,7,7,7,8,2,2,7,7,8,8,1),
	(1,1,1,8,7,14,14,7,14,14,7,7,7,7,9,7,14,9,14,7,8,9,7,7,7,7,7,7,9,8,14,1),
	(1,1,1,9,7,7,14,7,8,7,8,7,8,7,7,7,8,8,8,14,12,8,9,7,7,7,9,7,8,14,8,1),
	(1,1,1,7,7,8,9,7,8,9,14,14,8,8,9,8,8,9,14,14,12,8,8,7,14,9,8,7,7,7,8,1),
	(1,1,1,7,8,9,8,7,8,7,8,7,14,2,2,8,2,2,8,8,8,7,7,7,8,14,8,8,9,7,7,1),
	(1,1,1,7,9,7,7,7,7,7,9,14,8,7,7,7,7,7,8,9,7,7,12,7,7,8,2,2,8,9,7,1),
	(1,1,1,7,8,9,8,9,9,7,7,8,7,7,7,9,7,7,8,7,7,12,12,12,7,7,7,2,14,14,7,1),
	(1,1,1,7,7,8,8,9,9,7,7,7,7,8,8,8,8,7,8,14,7,7,12,7,7,14,7,2,14,7,7,1),
	(1,1,1,9,7,7,8,8,8,8,8,7,7,7,9,8,9,7,14,8,8,7,7,7,14,7,7,2,8,7,7,1),
	(1,1,1,9,9,7,8,8,8,7,9,8,9,7,7,8,8,7,7,7,8,8,7,14,2,2,7,8,9,9,9,1),
	(1,1,1,9,7,7,7,7,14,7,7,7,7,7,7,9,7,9,8,7,7,9,7,7,7,7,7,7,8,9,2,1),
	(1,1,1,7,7,8,12,7,14,14,14,12,8,9,7,7,7,7,9,7,7,7,9,8,7,2,9,7,9,2,2,1),
	(1,1,1,8,8,8,7,7,14,7,14,12,8,9,8,7,7,9,8,8,8,7,8,7,8,8,2,7,7,7,2,1),
	(1,1,1,8,8,7,7,9,8,7,8,12,8,8,7,7,8,9,9,8,7,7,7,7,12,8,2,2,8,7,8,1),
	(1,1,1,12,12,7,9,8,12,7,8,8,12,8,7,7,7,7,7,7,7,9,7,12,12,12,8,2,8,6,6,1),
	(1,1,1,12,12,7,7,7,7,7,7,12,12,8,8,9,8,12,12,12,12,8,8,12,12,12,8,2,8,6,6,1),
	(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1)
	);

constant nivel_2 : mem_matrix := (
	(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
	(1,1,1,9, 8, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 8, 7, 7, 7, 8, 7, 7, 7, 8, 7, 7, 7, 14,11,14,11,1),
	(1,1,1,9, 14,8, 14,14,7, 8, 7, 8, 7, 11,7, 7, 7, 8, 7, 14,9, 14,7, 7, 7, 14,7, 8, 2, 2, 2, 1),
	(1,1,1,9, 12,12,8, 7, 7, 14,7, 8, 14,8, 8, 8, 14,14,7, 8, 14,8, 7, 14,14,14,7, 8, 2, 8, 8, 1),
	(1,1,1,9, 14,14,8, 7, 14,7, 7, 8, 9, 9, 9, 14,9, 9, 7, 7, 7, 7, 7, 14,7, 14,7, 14,2, 11,11,1),
	(1,1,1,9, 8, 11,14,14,8, 8, 7, 9, 9, 14,9, 9, 9, 14,14,7, 8, 8, 8, 7, 7, 14,7, 8, 2, 8, 8, 1),
	(1,1,1,7, 7, 7, 7, 7, 7, 7, 7, 14,14,14,14,14,14,7, 14,7, 7, 7, 14,14,12,7, 7, 8, 7, 7, 7, 1),
	(1,1,1,7, 14,14,2, 14,14,14,7, 7, 7, 14,7, 7, 7, 7, 14,14,14,7, 14,7, 7, 7, 14,8, 14,8, 7, 1),
	(1,1,1,7, 14,11,11,14,2, 14,14,14,7, 14,7, 14,14,7, 7, 7, 7, 7, 14,14,12,7, 7, 7, 7, 8, 7, 1),
	(1,1,1,7, 14,11,11,14,7, 7, 7, 7, 7, 14,7, 7, 14,14,14,14,2, 9, 9, 2, 7, 11,14,8, 7, 8, 7, 1),
	(1,1,1,7, 14,11,11,14,7, 11,11,7, 14,14,14,7, 7, 7, 7, 7, 9, 11,11,9, 7, 14,7, 8, 7, 8, 7, 1),
	(1,1,1,7, 14,14,14,14,7, 7, 7, 7, 14,9, 9, 7, 14,7, 14,7, 9, 11,11,9, 7, 14,7, 8, 7, 7, 7, 1),
	(1,1,1,7, 14,2, 2, 7, 12,14,14,12,14,14,12,14,14,12,14,7, 2, 9, 9, 2, 7, 11,7, 8, 8, 8, 7, 1),
	(1,1,1,7, 14,14,14,7, 14,7, 7, 7, 7, 7, 7, 7, 9, 9, 7, 7, 8, 8, 7, 14,7, 14,7, 7, 7, 7, 7, 1),
	(1,1,1,7, 7, 7, 7, 7, 8, 7, 14,14,14,14,14,14,9, 8, 7, 14,7, 8, 7, 7, 7, 14,7, 8, 14,8, 8, 1),
	(1,1,1,8, 14,14,8, 7, 14,7, 14,7, 7, 7, 7, 7, 7, 14,12,8, 7, 14,8, 14,7, 11,7, 7, 7, 7, 7, 1),
	(1,1,1,7, 7, 7, 7, 7, 14,7, 7, 14,7, 8, 14,8, 14,14,14,14,7, 8, 7, 7, 7, 8, 14,14,8, 8, 7, 1),
	(1,1,1,7, 14,8, 14,14,8, 14,7, 14,7, 8, 7, 7, 7, 14,11,14,7, 8, 14,8, 7, 7, 7, 7, 7, 7, 7, 1),
	(1,1,1,7, 7, 7, 8, 7, 7, 7, 7, 14,7, 7, 7, 8, 7, 7, 2, 8, 7, 7, 7, 8, 14,8, 8, 14,8, 11,11,1),---
	(1,1,1,7, 8, 14,14,7, 14,14,14,14,14,14,14,14,14,14,7, 14,14,14,7, 14,7, 7, 7, 7, 14,9, 9, 1),
	(1,1,1,7, 7, 7, 7, 7, 7, 14,9, 9, 7, 7, 7, 7, 14,7, 7, 9, 11,14,7, 8, 7, 8, 14,7, 7, 7, 9, 1),
	(1,1,1,9, 14,9, 14,14,12,11,6, 6, 11,12,14,7, 14,7, 8, 14,14,14,7, 14,7, 14,7, 7, 14,8, 9, 1),
	(1,1,1,9, 14,12,12,14,12,11,6, 6, 11,12,14,7, 9, 7, 7, 7, 7, 7, 7, 7, 7, 14,7, 14,8, 9, 9, 1),
	(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1)
	);
	
constant nivel_3 : mem_matrix := (
	(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
	(1,1,1,7,7,7,8,7,7,7,7,7,7,7,7,12,12,12,7,7,7,7,7,7,7,12,7,7,7,7,12,1),
	(1,1,1,7,7,7,8,7,7,12,12,14,14,14,7,7,7,7,7,14,14,14,14,9,7,7,7,8,12,7,12,1),
	(1,1,1,9,7,8,12,7,7,12,14,14,2,2,8,8,8,8,8,2,2,2,2,8,8,8,8,7,7,7,7,1),
	(1,1,1,9,7,14,12,7,7,12,14,14,2,11,11,2,11,2,11,11,11,2,11,11,11,11,8,7,2,2,7,1),
	(1,1,1,7,7,14,12,7,7,12,12,14,2,11,7,7,7,7,7,7,7,7,7,7,7,7,8,7,2,2,7,1),
	(1,1,1,7,9,8,12,12,7,7,7,8,2,11,7,14,14,14,14,7,7,7,7,7,9,7,8,7,7,7,7,1),
	(1,1,1,7,9,11,8,12,12,12,7,8,2,11,7,7,7,7,7,7,9,9,9,7,7,7,8,7,7,7,7,1),
	(1,1,1,7,7,7,11,8,12,12,7,8,2,2,2,2,7,11,7,7,14,14,14,7,7,7,7,8,2,7,2,1),
	(1,1,1,9,7,7,11,8,11,11,7,8,2,2,2,2,7,7,7,7,7,7,7,7,11,11,7,7,8,7,7,1),
	(1,1,1,7,7,8,8,7,7,7,7,2,2,2,2,2,9,9,9,7,7,14,11,7,2,2,11,7,14,2,7,1),
	(1,1,1,7,8,7,7,7,11,7,7,2,2,2,2,2,6,6,9,7,7,14,11,7,2,2,11,7,14,7,7,1),
	(1,1,1,7,14,7,11,11,11,11,11,2,2,2,2,2,6,6,9,7,7,14,7,7,11,7,11,7,14,7,2,1),
	(1,1,1,7,8,7,7,7,7,7,7,8,2,2,2,2,9,9,9,7,7,14,7,7,11,7,7,7,8,7,2,1),
	(1,1,1,7,11,8,14,14,8,2,7,8,2,2,2,2,7,7,7,7,7,7,7,7,14,7,7,8,7,7,2,1),
	(1,1,1,7,7,7,7,7,7,8,7,7,8,8,2,2,7,7,7,2,7,7,2,7,14,7,8,2,7,2,2,1),
	(1,1,1,11,11,9,11,9,7,14,7,7,7,8,9,9,11,7,7,7,7,2,7,7,7,7,7,8,7,7,2,1),
	(1,1,1,11,11,11,7,7,7,8,7,2,7,2,8,9,14,8,2,7,7,7,7,7,2,7,7,7,8,7,7,1),
	(1,1,1,8,8,8,7,11,8,7,7,7,7,2,8,7,7,7,7,2,2,2,2,2,2,11,7,7,11,14,7,1),
	(1,1,1,12,7,7,7,11,8,12,2,2,7,2,8,7,9,9,7,7,7,7,7,7,7,7,11,7,11,14,7,1),
	(1,1,1,12,7,12,12,11,8,12,2,2,7,8,2,7,9,9,12,14,14,14,14,14,8,7,7,7,11,14,7,1),
	(1,1,1,12,7,12,12,2,2,7,7,7,7,8,2,7,7,7,7,2,11,11,9,9,8,8,8,8,8,8,7,1),
	(1,1,1,12,7,7,7,7,7,7,12,12,12,8,2,12,12,12,7,7,7,7,7,7,7,7,7,7,7,7,7,1),
	(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1)
	);
	
constant victoria : mem_matrix := (
	(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
	(1,1,1,1,11,12,12,12,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
	(1,1,1,11,12,12,12,12,12,12,12,12,1,11,12,12,1,1,11,12,12,12,1,1,11,12,11,12,1,1,1,1),
	(1,1,1,11,12,4,15,12,12,4,15,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1),
	(1,1,1,11,12,4,15,12,12,4,15,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1),
	(1,1,1,11,12,12,4,15,4,15,12,12,12,4,15,15,15,12,12,4,15,12,12,4,15,12,4,15,4,15,12,1),
	(1,1,1,11,12,12,4,15,4,15,12,12,4,15,12,12,4,15,12,4,15,12,12,4,15,12,12,12,12,12,12,1),
	(1,1,1,11,12,12,12,4,15,12,12,12,4,15,12,12,4,15,12,4,15,12,12,4,15,12,4,15,4,15,12,1),
	(1,1,1,11,12,12,12,4,15,12,12,12,4,15,12,12,4,15,12,4,15,12,12,4,15,12,12,4,15,12,12,1),
	(1,1,1,11,12,12,12,4,15,12,12,12,4,15,12,12,4,15,12,4,15,12,12,4,15,12,12,12,12,12,12,1),
	(1,1,1,11,12,12,12,4,15,12,12,12,12,4,15,15,15,12,12,12,4,15,15,15,12,12,12,12,12,12,1,1),
	(1,1,1,1,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1,1,1),
	(1,1,1,1,1,1,11,12,12,12,1,1,11,12,1,11,12,1,11,12,1,11,12,1,1,11,12,12,1,1,1,1),
	(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
	(1,1,1,1,11,12,12,12,12,12,12,12,1,11,12,12,1,11,12,12,1,11,12,12,1,11,12,12,12,1,1,1),
	(1,1,1,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1,1,1),
	(1,1,1,11,12,4,15,12,12,12,12,4,15,12,4,15,15,15,12,4,15,12,12,4,15,12,4,15,12,12,1,1),
	(1,1,1,11,12,4,15,12,4,15,12,4,15,12,12,4,15,12,12,4,15,15,12,4,15,12,4,15,12,12,12,1),
	(1,1,1,11,12,12,4,15,4,15,4,15,12,12,12,4,15,12,12,4,15,4,15,4,15,12,4,15,12,12,12,1),
	(1,1,1,11,12,12,4,15,4,15,4,15,12,12,12,4,15,12,12,4,15,12,4,15,15,12,12,12,12,12,12,1),
	(1,1,1,11,12,12,12,4,15,4,15,12,12,12,4,15,15,15,12,4,15,12,12,4,15,12,4,15,12,12,1,1),
	(1,1,1,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1,1,1),
	(1,1,1,1,11,12,12,12,1,11,12,12,1,11,12,1,11,12,1,11,12,1,11,12,12,1,11,12,1,1,1,1),
	(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1)
	);

constant game_over : mem_matrix := (
	(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
	(1,1,1,1,11,12,12,12,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
	(1,1,1,11,12,12,12,12,12,12,12,12,12,11,12,12,1,1,11,12,12,12,1,1,11,12,11,12,1,1,1,1),
	(1,1,1,11,12,2,15,15,15,15,15,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1),
	(1,1,1,11,12,2,15,12,12,2,15,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1),
	(1,1,1,11,12,2,15,12,12,12,12,12,12,2,15,15,12,12,12,2,15,2,15,12,12,12,2,15,15,12,12,1),
	(1,1,1,11,12,2,15,12,2,15,15,12,2,15,12,2,15,12,2,15,2,15,2,15,12,2,15,12,12,12,12,1),
	(1,1,1,11,12,2,15,12,12,2,15,12,2,15,15,15,15,12,2,15,2,15,2,15,12,2,15,15,12,12,12,1),
	(1,1,1,11,12,2,15,12,12,2,15,12,2,15,12,2,15,12,2,15,12,12,2,15,12,2,15,12,12,12,12,1),
	(1,1,1,11,12,2,15,15,15,15,15,12,2,15,12,2,15,12,2,15,12,12,2,15,12,12,2,15,15,12,12,1),
	(1,1,1,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1,1),
	(1,1,1,1,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1,1,1),
	(1,1,1,1,1,1,11,12,12,12,1,1,11,12,1,11,12,1,11,12,1,11,12,1,1,11,12,12,1,1,1,1),
	(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
	(1,1,1,1,11,12,12,12,12,12,12,12,1,11,12,12,1,11,12,12,1,11,12,12,1,11,12,12,12,1,1,1),
	(1,1,1,11,12,12,2,15,15,15,15,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1,1),
	(1,1,1,11,12,2,15,12,12,12,2,15,12,2,15,12,12,2,15,12,12,2,15,15,12,2,15,15,15,12,12,1),
	(1,1,1,11,12,2,15,12,12,12,2,15,12,2,15,12,12,2,15,12,2,15,12,12,12,2,15,12,2,15,12,1),
	(1,1,1,11,12,2,15,12,12,12,2,15,12,12,2,15,2,15,12,12,2,15,15,12,12,2,15,15,15,15,12,1),
	(1,1,1,11,12,2,15,12,12,12,2,15,12,12,2,15,2,15,12,12,2,15,12,12,12,2,15,12,2,15,12,1),
	(1,1,1,11,12,12,2,15,15,15,15,12,12,12,12,2,15,12,12,12,12,2,15,15,12,2,15,12,2,15,12,1),
	(1,1,1,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,1),
	(1,1,1,1,11,12,12,12,1,11,12,12,1,11,12,1,11,12,1,11,12,1,11,12,12,12,1,11,12,12,1,1),
	(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1)
	);

begin

	--Dependiendo del nivel se selecciona una de las memorias.
	process(NIVEL,FILA,COLUMNA)
	begin
		if(NIVEL = 0) then
			COLORES <= inicio(FILA,COLUMNA);
		elsif (NIVEL = 1) then
			COLORES <= nivel_1(FILA,COLUMNA);
		elsif (NIVEL = 2) then
			COLORES <= nivel_2(FILA,COLUMNA);
		elsif (NIVEL = 3) then
			COLORES <= nivel_3(FILA,COLUMNA);
		elsif (NIVEL = 4) then
			COLORES <= victoria(FILA,COLUMNA);
		else
			COLORES <= game_over(FILA,COLUMNA);
		end if;
	end process;

end Behavioral;

