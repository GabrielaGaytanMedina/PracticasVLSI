library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mem_prota is
    Port ( FILA  : in  integer;
           COLUMNA : in  integer;
           COLOR : out  integer);
end mem_prota;

architecture Behavioral of mem_prota is

type mem_matrix is array (0 to 31, 0 to 31) of integer;
constant memo : mem_matrix := (
	(0,0,0,0,0,0,0,5,5,5,5,5,5,5,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	(0,0,0,0,0,5,5,5,5,5,5,5,5,5,5,5,0,0,0,0,10,10,10,0,0,0,0,10,10,10,0,0),
	(0,0,0,0,5,5,5,5,5,5,5,5,5,5,5,5,5,0,10,10,10,10,10,10,0,0,10,10,10,10,10,0),
	(0,0,0,5,5,5,5,5,5,5,5,3,3,3,5,5,5,10,10,10,10,2,2,10,0,10,10,10,10,2,2,10),
	(0,0,5,5,5,3,3,3,5,5,5,5,3,3,5,5,5,10,10,10,10,2,1,10,10,10,10,10,10,2,1,10),
	(0,0,5,5,5,3,3,3,5,5,5,5,5,5,5,5,5,10,10,10,10,2,2,10,10,10,10,10,10,2,2,10),
	(0,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,10,10,10,10,10,10,0,10,10,10,10,10,10,10),
	(0,5,3,3,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,10,10,10,10,0,0,0,10,10,10,10,10,0),
	(5,5,3,5,5,5,2,2,2,5,5,5,5,5,5,5,5,5,5,5,13,13,10,0,0,0,0,10,13,13,13,0),
	(5,5,5,5,5,2,2,2,2,5,5,5,5,5,5,3,3,5,5,5,13,13,13,0,0,0,0,13,13,13,0,0),
	(5,5,5,5,2,2,2,2,2,2,2,5,5,5,5,5,3,3,5,5,5,13,13,13,0,0,0,13,13,13,0,0),
	(5,5,5,5,2,2,5,5,5,2,2,5,5,5,5,5,5,3,5,5,5,5,13,13,0,0,0,13,13,0,0,0),
	(5,5,5,5,2,2,5,5,5,5,2,2,5,5,5,5,5,5,5,5,5,5,13,13,0,0,0,13,13,0,0,0),
	(5,5,5,5,2,2,5,5,5,5,2,2,5,5,5,5,5,5,5,5,5,5,13,13,0,0,0,13,13,0,0,0),
	(5,5,5,5,2,2,5,5,5,5,5,2,2,5,5,5,5,5,5,5,5,5,13,13,0,0,0,13,13,0,0,0),
	(5,5,5,5,2,2,2,5,5,5,5,2,2,5,5,5,5,3,3,5,5,5,13,13,13,0,0,13,13,0,0,0),
	(5,5,5,5,5,2,2,2,5,5,5,2,2,5,5,5,5,3,3,5,5,5,0,13,13,0,0,13,13,0,0,0),
	(5,5,5,5,5,5,2,2,5,5,5,2,2,5,5,5,5,5,5,5,5,5,0,13,13,0,0,13,13,0,0,0),
	(5,5,5,5,5,5,5,5,5,5,5,2,2,2,5,5,5,5,5,5,5,5,0,13,13,0,0,13,13,0,0,0),
	(0,5,5,5,5,5,5,5,5,5,5,5,2,2,5,5,5,5,5,5,5,5,0,13,13,0,0,13,13,0,0,0),
	(0,5,5,5,5,5,5,5,5,5,5,5,2,2,5,5,5,5,5,5,5,5,0,13,13,0,0,13,13,0,0,0),
	(0,5,5,5,5,5,5,5,5,5,5,5,2,2,5,5,5,5,5,5,5,5,0,13,13,0,0,13,13,0,0,0),
	(0,0,5,5,5,5,5,5,5,5,5,5,2,2,5,5,5,5,5,5,5,0,0,13,13,0,0,13,13,0,0,0),
	(0,0,5,5,5,5,5,5,5,5,5,5,2,2,5,5,5,5,5,5,5,0,0,13,13,0,13,13,0,0,0,0),
	(0,0,0,5,5,5,5,5,5,5,5,5,2,2,5,5,5,5,5,5,0,0,0,13,13,0,13,13,0,0,0,0),
	(0,0,0,0,5,5,5,5,5,5,5,5,2,2,5,5,5,5,5,5,0,0,0,13,13,0,13,13,0,0,0,0),
	(0,0,0,0,5,5,5,5,5,5,5,2,2,5,5,5,5,5,5,0,0,0,0,13,13,0,13,13,0,0,0,0),
	(0,0,0,0,0,5,5,5,5,5,2,2,2,5,5,5,5,13,13,13,13,13,13,13,13,0,13,13,0,0,0,0),
	(10,10,10,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,0,0),
	(10,10,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,10,0,0),
	(0,10,10,13,13,13,13,10,10,13,13,13,13,10,13,13,13,13,10,10,13,13,13,10,10,13,13,13,13,13,10,0),
	(0,0,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10)
	);

begin

	COLOR <= memo(FILA,COLUMNA);

end Behavioral;

